.title KiCad schematic
.include "C:/AE/TLP291-4/TLP291_4.mod"
.include "C:/AE/TLP291-4/ceu4j2x7r1h104m125ae_p.mod"
.include "C:/AE/TLP291-4/lmx24_lm2902.lib"
XU3 /LIN /DV2 VCC 0 /OA2 LMX24_LM2902
R6 /DV1 /DV2 {RDIV2}
XU2 /LIN /DV1 VCC 0 /OA1 LMX24_LM2902
R2 /K2 /OA2 {RK}
R1 /K1 /OA1 {RK}
R5 VCC /DV1 {RDIV1}
R8 /DV3 /DV4 {RDIV4}
R7 /DV2 /DV3 {RDIV3}
R3 /K3 /OA3 {RK}
XU5 /LIN /DV4 VCC 0 /OA4 LMX24_LM2902
XU4 /LIN /DV3 VCC 0 /OA3 LMX24_LM2902
R4 /K4 /OA4 {RK}
R9 /DV4 0 {RDIV5}
R12 VCC /LEXT {RPOWER}
R10 /LIN 0 {RREF}
R11 /LIN /LEXT {RSER}
XU6 /LIN 0 CEU4J2X7R1H104M125AE_p
R13 /LEXT 0 {RSTATE}
XU1 VCC /K1 VCC /K2 VCC /K3 VCC /K4 0 /OPT4 0 /OPT3 0 /OPT2 0 /OPT1 TLP291_4
R14 VDC /OPT1 {RPU}
R17 VDC /OPT4 {RPU}
R16 VDC /OPT3 {RPU}
R15 VDC /OPT2 {RPU}
XU7 VCC 0 CEU4J2X7R1H104M125AE_p
V1 VCC 0 DC {VSOURCE}
V2 VDC 0 DC {VDIG}
.end
